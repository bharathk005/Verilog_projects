`timescale 1ns / 1ps

module tester1_1();

endmodule
