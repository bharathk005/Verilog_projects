`timescale 1ns / 1ps

module tester1();

endmodule