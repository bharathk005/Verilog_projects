`timescale 1ns / 1ps

module mult(a,b,c,d);
input [0:15] a;
input [0:15] b;
input c;
output reg [0:15]d;

reg [0:15] r1;
reg [0:15] r3;
reg [0:15] r2;
reg [0:15] r22;
always@(*)
begin
/*	r1 <= a[3:15]*b[3:15];
	r2 <= ((a[0:2]*b[3:15])+(b[0:2]*a[3:15]))/10;
	r22 <= (a[0:2]*b[3:15])+(b[0:2]*a[3:15])-((((a[0:2]*b[3:15])+(b[0:2]*a[3:15]))/10)*10);
	r3 <= a[0:2]*b[0:2];
*/
	d[0:2] <= (a[0:2]*b[0:2])+(a[0:2]*b[3:15])+(b[0:2]*a[3:15])-((((a[0:2]*b[3:15])+(b[0:2]*a[3:15]))/10)*10);
	d[3:15] <= (a[3:15]*b[3:15])+(((a[0:2]*b[3:15])+(b[0:2]*a[3:15]))/10);
end	
//assign d[0:2] = r3+r22;
//assign d[3:15] = r1+r2;
endmodule
