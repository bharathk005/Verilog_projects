`timescale 1ns / 1ps

module vControl(
    );


endmodule
